`include "player1.v"
module finiteStateMachine (
    input health1,
    input health2,
    input clk,
    input action1,
    input action2
);
player1,

endmodule