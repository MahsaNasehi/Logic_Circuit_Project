`include "player1"
module finiteStateMachine (
    input health1,
    input health2,
    input clk,
    input action1,
    input action2
);

endmodule